library verilog;
use verilog.vl_types.all;
entity mux_21_vlg_vec_tst is
end mux_21_vlg_vec_tst;
