library verilog;
use verilog.vl_types.all;
entity Final_vlg_check_tst is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        DIG0            : in     vl_logic;
        DIG1            : in     vl_logic;
        DIG2            : in     vl_logic;
        DIG3            : in     vl_logic;
        e               : in     vl_logic;
        f               : in     vl_logic;
        g               : in     vl_logic;
        LED0            : in     vl_logic;
        LED1            : in     vl_logic;
        LED2            : in     vl_logic;
        LED3            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Final_vlg_check_tst;
