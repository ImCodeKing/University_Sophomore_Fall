library verilog;
use verilog.vl_types.all;
entity Final_vlg_vec_tst is
end Final_vlg_vec_tst;
