library verilog;
use verilog.vl_types.all;
entity mux_21_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux_21_vlg_check_tst;
