library verilog;
use verilog.vl_types.all;
entity AddAndMinus_vlg_tst is
end AddAndMinus_vlg_tst;
