library verilog;
use verilog.vl_types.all;
entity AddAndMinus_vlg_vec_tst is
end AddAndMinus_vlg_vec_tst;
